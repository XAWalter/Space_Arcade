`timescale 1ns/1ps
module uart_rx_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, uart_rx_tb);
	end
endmodule

