`timescale 1ns/1ps
module bt_control_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, bt_control_tb);
	end
endmodule

