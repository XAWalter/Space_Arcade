`timescale 1ns/1ps
module audio_control_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, audio_control_tb);
	end
endmodule

