`timescale 1ns/1ps
module spi_interface_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, spi_interface_tb);
	end
endmodule

