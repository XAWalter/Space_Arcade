`timescale 1ns/1ps
module clock_divider_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, clock_divider_tb);
	end
endmodule

